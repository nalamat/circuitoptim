Sample Optimization of RLC circuit
vs  vs  gnd ac  1
r1  out gnd 1k
l1  a   out 162u
c1  vs  a   752u
.ac lin 3k  1  5k
.option post = 1
.end