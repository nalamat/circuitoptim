Sample circuit of series RLC
vs  vs  gnd ac  1
r1  out gnd [10]     ** [1      1meg    dec]
l1  a   out [1m]     ** [1u     10m     dec]
c1  vs  a   [10u]    ** [10p    100u    lin]
.ac lin 3k  1  5k
.end