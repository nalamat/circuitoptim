Sample circuit of series RLC
vs  vs  gnd ac  1
r1  out gnd [10]     ** [1      1e6    dec]
l1  a   out [1e-3]   ** [1e-6   10e-3  dec]
c1  vs  a   [10e-6]  ** [10e-12 100e-6 dec]
.ac lin 3k  1  5k
.end